module led_blink (
    input clk,          // 50MHz onboard clock
    output reg led1,    // LED1 output
    output reg led2,    // LED2 output
    output reg led3     // LED3 output
);

// Clock divider for 0.5s intervals (50MHz → 1Hz enable)
reg [24:0] counter;
wire enable = (counter == 25'd24_999_999);  // 0.5s at 50MHz

// 2-bit state register for LED control
reg [1:0] state;

always @(posedge clk) begin
    // Clock divider logic
    counter <= (enable) ? 0 : counter + 1;
    
    // State machine
    if(enable) begin
        state <= (state == 2'b10) ? 2'b00 : state + 1;
    end
end

// LED output logic
always @(*) begin
    case(state)
        2'b00: {led1, led2, led3} = 3'b100;  // LED1 on
        2'b01: {led1, led2, led3} = 3'b010;  // LED2 on
        2'b10: {led1, led2, led3} = 3'b001;  // LED3 on
        default: {led1, led2, led3} = 3'b000; // All off
    endcase
end

endmodule